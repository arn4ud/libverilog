module test0
endmodule