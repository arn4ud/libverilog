module test1(input i0, input i1, output O);
endmodule