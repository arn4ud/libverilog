module test1(i0, i1, O);
input i0;
input i1;
input O;

endmodule